configuration NZPsplit_config of NZPsplit is
   for untitled
   end for;
end NZPsplit_config;