configuration StoreMux_config of StoreMux is
   for untitled
   end for;
end StoreMux_config;