configuration Plus2_config of Plus2 is
   for untitled
   end for;
end Plus2_config;