configuration Reg16_config of Reg16 is
   for untitled
   end for;
end Reg16_config;