--
-- VHDL Architecture ece411.SEXT11.untitled
--
-- Created:
--          by - wheele11.ews (gelib-057-06.ews.illinois.edu)
--          at - 20:48:31 03/09/12
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY SEXT11 IS
   PORT( 
      in11   : IN     std_logic_vector (10 DOWNTO 0);
      output : OUT    LC3b_word
   );

-- Declarations

END SEXT11 ;

--
-- VHDL Architecture ece411.SEXT11.struct
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

LIBRARY mp3lib;

ARCHITECTURE struct OF SEXT11 IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL one  : STD_LOGIC;
   SIGNAL zero : STD_LOGIC;


   -- Component Declarations
   COMPONENT TRISTATE1_H
   PORT (
      A  : IN     STD_LOGIC ;
      EN : IN     STD_LOGIC ;
      F  : OUT    STD_LOGIC 
   );
   END COMPONENT;
   COMPONENT TRISTATE1_L
   PORT (
      A  : IN     STD_LOGIC ;
      EN : IN     STD_LOGIC ;
      F  : OUT    STD_LOGIC 
   );
   END COMPONENT;


BEGIN
   -- Architecture concurrent statements
   -- HDL Embedded Text Block 2 eb2
   output(11 downto 0) <= in11 & '0';
   zero <= '0';
   one  <= '1';


   -- Instance port mappings.

   g3: FOR i IN 12 TO 15 GENERATE
   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : TRISTATE1_H USE ENTITY mp3lib.TRISTATE1_H;
   -- pragma synthesis_on

   BEGIN
      U_3 : TRISTATE1_H
         PORT MAP (
            A  => one,
            EN => in11(10),
            F  => output(i)
         );
   END GENERATE g3;

   g4: FOR i IN 12 TO 15 GENERATE
   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : TRISTATE1_L USE ENTITY mp3lib.TRISTATE1_L;
   -- pragma synthesis_on

   BEGIN
      U_0 : TRISTATE1_L
         PORT MAP (
            A  => zero,
            EN => in11(10),
            F  => output(i)
         );
   END GENERATE g4;

END struct;
