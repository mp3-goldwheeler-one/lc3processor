configuration GenCC_config of GenCC is
   for untitled
   end for;
end GenCC_config;