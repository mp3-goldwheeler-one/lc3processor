--
-- VHDL Architecture ece411.Memory.untitled
--
-- Created:
--          by - goldste6.UNKNOWN (linux4.ews.illinois.edu)
--          at - 20:21:18 01/18/12
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Memory IS
   PORT( 
      CLK              : IN     std_logic;
      RESET_L          : IN     STD_LOGIC;
      data_mread_l     : IN     std_logic;
      data_mwrite_l    : IN     STD_LOGIC;
      data_pm_addr     : IN     LC3B_WORD;
      data_pm_dataout  : IN     LC3B_OWORD;
      instr_mread_l    : IN     std_logic;
      instr_mwrite_l   : IN     STD_LOGIC;
      instr_pm_addr    : IN     LC3b_word;
      instr_pm_dataout : IN     lc3b_oword;
      data_in          : OUT    LC3B_OWORD;
      data_resp_h      : OUT    std_logic;
      instr_in         : OUT    LC3B_OWORD;
      instr_resp_h     : OUT    std_logic
   );

-- Declarations

END Memory ;

--
-- VHDL Architecture ece411.Memory.struct
--
-- Created:
--          by - one1.ews (gelib-057-16.ews.illinois.edu)
--          at - 17:57:47 04/26/12
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

LIBRARY ece411;
LIBRARY mp3lib;

ARCHITECTURE struct OF Memory IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL ADDRESS        : LC3B_WORD;
   SIGNAL DATAIN         : LC3B_OWORD;
   SIGNAL DATAOUT        : LC3B_OWORD;
   SIGNAL D_PMADDRESS    : LC3B_WORD;
   SIGNAL D_PMDATAOUT    : LC3B_OWORD;
   SIGNAL D_PMREAD_L     : std_logic;
   SIGNAL D_PMRESP_H     : std_logic;
   SIGNAL D_PMWRITE_L    : std_logic;
   SIGNAL FIXED_PMRESP_H : STD_LOGIC;
   SIGNAL I_PMADDRESS    : LC3B_WORD;
   SIGNAL I_PMDATAOUT    : LC3B_OWORD;
   SIGNAL I_PMREAD_L     : std_logic;
   SIGNAL I_PMRESP_H     : STD_LOGIC;
   SIGNAL I_PMWRITE_L    : std_logic;
   SIGNAL MREAD_L        : STD_LOGIC;
   SIGNAL MRESP_H        : STD_LOGIC;
   SIGNAL MWRITE_L       : STD_LOGIC;
   SIGNAL PMADDRESS      : LC3B_WORD;
   SIGNAL PMDATAIN       : LC3B_PWORD;
   SIGNAL PMDATAOUT      : LC3B_PWORD;
   SIGNAL PMREAD_L       : STD_LOGIC;
   SIGNAL PMRESP_H       : std_logic;
   SIGNAL PMWRITE_L      : STD_LOGIC;


   -- Component Declarations
   COMPONENT Cache_Arbiter
   PORT (
      CLK         : IN     std_logic ;
      D_PMADDRESS : IN     LC3B_WORD ;
      D_PMDATAOUT : IN     LC3B_OWORD ;
      D_PMREAD_L  : IN     std_logic ;
      D_PMWRITE_L : IN     std_logic ;
      I_PMADDRESS : IN     LC3B_WORD ;
      I_PMDATAOUT : IN     LC3B_OWORD ;
      I_PMREAD_L  : IN     std_logic ;
      I_PMWRITE_L : IN     std_logic ;
      MRESP_H     : IN     STD_LOGIC ;
      RESET_L     : IN     STD_LOGIC ;
      ADDRESS     : OUT    LC3B_WORD ;
      DATAOUT     : OUT    LC3B_OWORD ;
      D_PMRESP_H  : OUT    std_logic ;
      I_PMRESP_H  : OUT    STD_LOGIC ;
      MREAD_L     : OUT    STD_LOGIC ;
      MWRITE_L    : OUT    STD_LOGIC 
   );
   END COMPONENT;
   COMPONENT Fix_pmresp_h
   PORT (
      PMRESP_H       : IN     std_logic ;
      FIXED_PMRESP_H : OUT    STD_LOGIC 
   );
   END COMPONENT;
   COMPONENT L2_Cache
   PORT (
      ADDRESS   : IN     LC3B_WORD ;
      CLK       : IN     std_logic ;
      Dataout   : IN     LC3B_OWORD ;
      MREAD_L   : IN     std_logic ;
      MWRITE_L  : IN     std_logic ;
      PMDATAIN  : IN     LC3B_PWORD ;
      PMRESP_H  : IN     std_logic ;
      RESET_L   : IN     std_logic ;
      DATAIN    : OUT    LC3B_OWORD ;
      MRESP_H   : OUT    std_logic ;
      PMADDRESS : OUT    LC3B_WORD ;
      PMDATAOUT : OUT    LC3B_PWORD ;
      PMREAD_L  : OUT    std_logic ;
      PMWRITE_L : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT DRAM256
   PORT (
      ADDRESS  : IN     LC3B_WORD ;
      DATAOUT  : IN     LC3B_PWORD ;
      MREAD_L  : IN     STD_LOGIC ;
      MWRITE_L : IN     STD_LOGIC ;
      RESET_L  : IN     STD_LOGIC ;
      DATAIN   : OUT    LC3B_PWORD ;
      MRESP_H  : OUT    STD_LOGIC 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Cache_Arbiter USE ENTITY ece411.Cache_Arbiter;
   FOR ALL : DRAM256 USE ENTITY mp3lib.DRAM256;
   FOR ALL : Fix_pmresp_h USE ENTITY ece411.Fix_pmresp_h;
   FOR ALL : L2_Cache USE ENTITY ece411.L2_Cache;
   -- pragma synthesis_on


BEGIN
   -- Architecture concurrent statements
   -- HDL Embedded Text Block 1 eb1
   I_PMREAD_L    <= instr_mread_l;
   I_PMWRITE_L   <= instr_mwrite_l;
   I_PMADDRESS   <= instr_pm_addr;
   I_PMDATAOUT   <= instr_pm_dataout;
   instr_in      <= DATAIN;
   instr_resp_h  <= I_PMRESP_H;

   -- HDL Embedded Text Block 2 eb2
   D_PMREAD_L   <= data_mread_l;
   D_PMWRITE_L  <= data_mwrite_l;
   D_PMADDRESS  <= data_pm_addr;
   D_PMDATAOUT  <= data_pm_dataout;
   data_in      <= DATAIN;
   data_resp_h  <= D_PMRESP_H;


   -- Instance port mappings.
   arbiter : Cache_Arbiter
      PORT MAP (
         CLK         => CLK,
         D_PMADDRESS => D_PMADDRESS,
         D_PMDATAOUT => D_PMDATAOUT,
         D_PMREAD_L  => D_PMREAD_L,
         D_PMWRITE_L => D_PMWRITE_L,
         I_PMADDRESS => I_PMADDRESS,
         I_PMDATAOUT => I_PMDATAOUT,
         I_PMREAD_L  => I_PMREAD_L,
         I_PMWRITE_L => I_PMWRITE_L,
         MRESP_H     => MRESP_H,
         RESET_L     => RESET_L,
         ADDRESS     => ADDRESS,
         DATAOUT     => DATAOUT,
         D_PMRESP_H  => D_PMRESP_H,
         I_PMRESP_H  => I_PMRESP_H,
         MREAD_L     => MREAD_L,
         MWRITE_L    => MWRITE_L
      );
   fixResponse : Fix_pmresp_h
      PORT MAP (
         PMRESP_H       => PMRESP_H,
         FIXED_PMRESP_H => FIXED_PMRESP_H
      );
   l2 : L2_Cache
      PORT MAP (
         ADDRESS   => ADDRESS,
         CLK       => CLK,
         Dataout   => DATAOUT,
         MREAD_L   => MREAD_L,
         MWRITE_L  => MWRITE_L,
         PMDATAIN  => PMDATAIN,
         PMRESP_H  => FIXED_PMRESP_H,
         RESET_L   => RESET_L,
         DATAIN    => DATAIN,
         MRESP_H   => MRESP_H,
         PMADDRESS => PMADDRESS,
         PMDATAOUT => PMDATAOUT,
         PMREAD_L  => PMREAD_L,
         PMWRITE_L => PMWRITE_L
      );
   Phys_Mem : DRAM256
      PORT MAP (
         ADDRESS  => PMADDRESS,
         DATAOUT  => PMDATAOUT,
         MREAD_L  => PMREAD_L,
         MWRITE_L => PMWRITE_L,
         RESET_L  => RESET_L,
         DATAIN   => PMDATAIN,
         MRESP_H  => PMRESP_H
      );

END struct;
