
--
ARCHITECTURE untitled OF Cache_Datapath IS
BEGIN
END ARCHITECTURE untitled;

