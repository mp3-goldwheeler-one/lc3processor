
--
ARCHITECTURE untitled OF BTB_Datapath IS
BEGIN
END ARCHITECTURE untitled;

