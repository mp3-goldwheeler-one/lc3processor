configuration ADJ6_config of ADJ6 is
   for untitled
   end for;
end ADJ6_config;