--
-- VHDL Architecture ece411.SEXT9.untitled
--
-- Created:
--          by - wheele11.ews (gelib-057-06.ews.illinois.edu)
--          at - 20:44:12 03/09/12
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY SEXT9 IS
   PORT( 
      in9    : IN     std_logic_vector (8 DOWNTO 0);
      output : OUT    std_logic_vector (15 DOWNTO 0)
   );

-- Declarations

END SEXT9 ;

--
-- VHDL Architecture ece411.SEXT9.struct
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

LIBRARY mp3lib;

ARCHITECTURE struct OF SEXT9 IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL one  : STD_LOGIC;
   SIGNAL zero : STD_LOGIC;


   -- Component Declarations
   COMPONENT TRISTATE1_H
   PORT (
      A  : IN     STD_LOGIC ;
      EN : IN     STD_LOGIC ;
      F  : OUT    STD_LOGIC 
   );
   END COMPONENT;
   COMPONENT TRISTATE1_L
   PORT (
      A  : IN     STD_LOGIC ;
      EN : IN     STD_LOGIC ;
      F  : OUT    STD_LOGIC 
   );
   END COMPONENT;


BEGIN
   -- Architecture concurrent statements
   -- HDL Embedded Text Block 1 eb1
   output(9 downto 0) <= in9 & '0';
   zero <= '0';
   one <= '1';


   -- Instance port mappings.

   g2: FOR i IN 10 TO 15 GENERATE
   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : TRISTATE1_H USE ENTITY mp3lib.TRISTATE1_H;
   -- pragma synthesis_on

   BEGIN
      U_3 : TRISTATE1_H
         PORT MAP (
            A  => one,
            EN => in9(8),
            F  => output(i)
         );
   END GENERATE g2;

   g3: FOR i IN 10 TO 15 GENERATE
   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : TRISTATE1_L USE ENTITY mp3lib.TRISTATE1_L;
   -- pragma synthesis_on

   BEGIN
      U_0 : TRISTATE1_L
         PORT MAP (
            A  => zero,
            EN => in9(8),
            F  => output(i)
         );
   END GENERATE g3;

END struct;
