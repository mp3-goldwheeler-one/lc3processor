--
-- VHDL Architecture ece411.id_reg_pipe.untitled
--
-- Created:
--          by - wheele11.ews (gelib-057-17.ews.illinois.edu)
--          at - 22:42:41 02/29/12
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY decode_exec_pipe IS
   PORT( 
      CLK                   : IN     std_logic;
      RESET_L               : IN     STD_LOGIC;
      decode_alumux_sel     : IN     STD_LOGIC_VECTOR (1 DOWNTO 0);
      decode_aluop          : IN     LC3b_aluop;
      decode_dr             : IN     LC3B_REG;
      decode_instr          : IN     STD_LOGIC_VECTOR (15 DOWNTO 0);
      decode_load_jump_pc   : IN     STD_LOGIC;
      decode_opcode         : IN     LC3b_opcode;
      decode_pc             : IN     LC3b_word;
      decode_read           : IN     std_logic;
      decode_regwrite       : IN     std_logic;
      decode_set_cc         : IN     std_logic;
      decode_shift_imm      : IN     STD_LOGIC;
      decode_src_a          : IN     LC3b_word;
      decode_src_b          : IN     LC3b_word;
      decode_use_offset11   : IN     STD_LOGIC;
      decode_use_pc_adder   : IN     STD_LOGIC;
      decode_write_byte     : IN     std_logic;
      decode_write_word     : IN     std_logic;
      load_decode_exec_pipe : IN     STD_LOGIC;
      exec_alumux_sel       : OUT    LC3b_4mux_sel;
      exec_aluop            : OUT    LC3B_ALUOP;
      exec_dr               : OUT    LC3B_REG;
      exec_instr            : OUT    LC3b_word;
      exec_load_jump_pc     : OUT    STD_LOGIC;
      exec_opcode           : OUT    LC3b_opcode;
      exec_pc               : OUT    LC3b_word;
      exec_read             : OUT    std_logic;
      exec_regwrite         : OUT    STD_LOGIC;
      exec_set_cc           : OUT    std_logic;
      exec_shift_imm        : OUT    STD_LOGIC;
      exec_src_a            : OUT    LC3b_word;
      exec_src_b            : OUT    LC3b_word;
      exec_use_offset11     : OUT    std_logic;
      exec_use_pc_adder     : OUT    std_logic;
      exec_write_byte       : OUT    std_logic;
      exec_write_word       : OUT    std_logic
   );

-- Declarations

END decode_exec_pipe ;

--
-- VHDL Architecture ece411.decode_exec_pipe.struct
--
-- Created:
--          by - goldste6.ews (gelib-057-26.ews.illinois.edu)
--          at - 19:47:43 03/13/12
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

LIBRARY mp3lib;

ARCHITECTURE struct OF decode_exec_pipe IS

   -- Architecture declarations

   -- Internal signal declarations


   -- Component Declarations
   COMPONENT REG1
   PORT (
      RESET_L : IN     STD_LOGIC ;
      A       : IN     STD_LOGIC ;
      EN      : IN     STD_LOGIC ;
      CLK     : IN     STD_LOGIC ;
      F       : OUT    STD_LOGIC 
   );
   END COMPONENT;
   COMPONENT REG16
   PORT (
      RESET_L : IN     STD_LOGIC ;
      A       : IN     STD_LOGIC_VECTOR (15 DOWNTO 0);
      EN      : IN     STD_LOGIC ;
      CLK     : IN     STD_LOGIC ;
      F       : OUT    STD_LOGIC_VECTOR (15 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT REG2
   PORT (
      RESET_L : IN     STD_LOGIC ;
      A       : IN     STD_LOGIC_VECTOR (1 DOWNTO 0);
      EN      : IN     STD_LOGIC ;
      CLK     : IN     STD_LOGIC ;
      F       : OUT    STD_LOGIC_VECTOR (1 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT REG3
   PORT (
      RESET_L : IN     STD_LOGIC ;
      A       : IN     STD_LOGIC_VECTOR (2 DOWNTO 0);
      EN      : IN     STD_LOGIC ;
      CLK     : IN     STD_LOGIC ;
      F       : OUT    STD_LOGIC_VECTOR (2 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT REG4
   PORT (
      RESET_L : IN     STD_LOGIC ;
      A       : IN     STD_LOGIC_VECTOR (3 DOWNTO 0);
      EN      : IN     STD_LOGIC ;
      CLK     : IN     STD_LOGIC ;
      F       : OUT    STD_LOGIC_VECTOR (3 DOWNTO 0)
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : REG1 USE ENTITY mp3lib.REG1;
   FOR ALL : REG16 USE ENTITY mp3lib.REG16;
   FOR ALL : REG2 USE ENTITY mp3lib.REG2;
   FOR ALL : REG3 USE ENTITY mp3lib.REG3;
   FOR ALL : REG4 USE ENTITY mp3lib.REG4;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   U_5 : REG1
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_regwrite,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_regwrite
      );
   U_9 : REG1
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_shift_imm,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_shift_imm
      );
   U_11 : REG1
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_use_offset11,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_use_offset11
      );
   U_12 : REG1
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_use_pc_adder,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_use_pc_adder
      );
   U_13 : REG1
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_load_jump_pc,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_load_jump_pc
      );
   U_14 : REG1
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_set_cc,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_set_cc
      );
   U_15 : REG1
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_write_byte,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_write_byte
      );
   U_17 : REG1
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_read,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_read
      );
   U_18 : REG1
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_write_word,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_write_word
      );
   U_0 : REG16
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_src_a,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_src_a
      );
   U_1 : REG16
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_src_b,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_src_b
      );
   U_2 : REG16
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_pc,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_pc
      );
   U_3 : REG16
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_instr,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_instr
      );
   U_10 : REG2
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_alumux_sel,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_alumux_sel
      );
   U_6 : REG3
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_aluop,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_aluop
      );
   U_7 : REG3
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_dr,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_dr
      );
   U_4 : REG4
      PORT MAP (
         RESET_L => RESET_L,
         A       => decode_opcode,
         EN      => load_decode_exec_pipe,
         CLK     => CLK,
         F       => exec_opcode
      );

END struct;
