configuration RegFile_config of RegFile is
   for untitled
   end for;
end RegFile_config;