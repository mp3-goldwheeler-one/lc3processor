configuration WordMux2_config of WordMux2 is
   for untitled
   end for;
end WordMux2_config;