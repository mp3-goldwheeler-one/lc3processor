configuration ALU_config of ALU is
   for untitled
   end for;
end ALU_config;