configuration ADJ9_config of ADJ9 is
   for untitled
   end for;
end ADJ9_config;