--
-- VHDL Architecture ece411.GenCC.untitled
--
-- Created:
--          by - goldste6.UNKNOWN (linux4.ews.illinois.edu)
--          at - 20:35:10 01/18/12
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY GenCC IS
   PORT( 
      WordIn  : IN     LC3b_word;
      nzp     : OUT    LC3b_cc
   );

-- Declarations

END GenCC ;

--
-- VHDL Architecture ece411.GenCC.struct
--
-- Created:
--          by - goldste6.ews (linux5.ews.illinois.edu)
--          at - 22:30:30 04/06/12
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

LIBRARY mp3lib;

ARCHITECTURE struct OF GenCC IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL zero_16 : LC3B_WORD;
   SIGNAL z       : STD_LOGIC;
   SIGNAL n       : STD_LOGIC;
   SIGNAL p       : STD_LOGIC;


   -- Component Declarations
   COMPONENT COMP16
   PORT (
      A : IN     LC3B_WORD ;
      B : IN     LC3B_WORD ;
      F : OUT    STD_LOGIC 
   );
   END COMPONENT;
   COMPONENT NOR2
   PORT (
      A : IN     STD_LOGIC ;
      B : IN     STD_LOGIC ;
      F : OUT    STD_LOGIC 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : COMP16 USE ENTITY mp3lib.COMP16;
   FOR ALL : NOR2 USE ENTITY mp3lib.NOR2;
   -- pragma synthesis_on


BEGIN
   -- Architecture concurrent statements
   -- HDL Embedded Text Block 1 eb1
   -- n and nzp generation
   n <= WordIn(15);
   nzp <= n & z & p;
   zero_16 <= x"0000";           


   -- Instance port mappings.
   U_1 : COMP16
      PORT MAP (
         A => WordIn,
         B => zero_16,
         F => z
      );
   U_0 : NOR2
      PORT MAP (
         A => z,
         B => n,
         F => p
      );

END struct;
