configuration BRadd_config of BRadd is
   for untitled
   end for;
end BRadd_config;