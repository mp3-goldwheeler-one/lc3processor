--
-- VHDL Architecture ece411.Memory.untitled
--
-- Created:
--          by - goldste6.UNKNOWN (linux4.ews.illinois.edu)
--          at - 20:21:18 01/18/12
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Memory IS
   PORT( 
      CLK             : IN     std_logic;
      Dataout         : IN     LC3b_word;
      RESET_L         : IN     STD_LOGIC;
      data_addr       : IN     LC3b_word;
      data_mread_l    : IN     std_logic;
      data_mwriteh_l  : IN     std_logic;
      data_mwritel_l  : IN     std_logic;
      instr_addr      : IN     LC3b_word;
      instr_mread_l   : IN     std_logic;
      instr_mwriteh_l : IN     std_logic;
      instr_mwritel_l : IN     std_logic;
      instr_out       : IN     std_logic;
      DATAIN          : OUT    std_logic;
      data_resp_h     : OUT    std_logic;
      instr_in        : OUT    LC3B_WORD;
      instr_resp_h    : OUT    std_logic
   );

-- Declarations

END Memory ;

--
-- VHDL Architecture ece411.Memory.struct
--
-- Created:
--          by - wheele11.ews (gelib-057-18.ews.illinois.edu)
--          at - 23:36:24 03/07/12
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

LIBRARY ece411;

ARCHITECTURE struct OF Memory IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL Address         : LC3b_word;
   SIGNAL DATAIN_internal : LC3b_word;
   SIGNAL Dirty           : std_logic;
   SIGNAL MREAD_L         : std_logic;
   SIGNAL MRESP_H         : std_logic;
   SIGNAL MWRITEH_L       : std_logic;
   SIGNAL MWRITEL_L       : std_logic;
   SIGNAL PMADDRESS       : LC3B_WORD;
   SIGNAL PMDATAIN        : LC3B_OWORD;
   SIGNAL PMDATAOUT       : LC3B_OWORD;
   SIGNAL PMREAD_L        : STD_LOGIC;
   SIGNAL PMRESP_H        : STD_LOGIC;
   SIGNAL PMWRITE_L       : STD_LOGIC;
   SIGNAL in_idlehit      : std_logic;
   SIGNAL in_load         : std_logic;
   SIGNAL in_writeback    : std_logic;
   SIGNAL miss            : std_logic;


   -- Component Declarations
   COMPONENT Cache_Controller
   PORT (
      CLK          : IN     std_logic ;
      Dirty        : IN     std_logic ;
      PMRESP_H     : IN     STD_LOGIC ;
      RESET_L      : IN     STD_LOGIC ;
      miss         : IN     std_logic ;
      PMREAD_L     : OUT    STD_LOGIC ;
      PMWRITE_L    : OUT    STD_LOGIC ;
      in_idlehit   : OUT    std_logic ;
      in_load      : OUT    std_logic ;
      in_writeback : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Cache_Datapath
   PORT (
      Address         : IN     LC3b_word ;
      CLK             : IN     std_logic ;
      Dataout         : IN     LC3b_word ;
      MREAD_L         : IN     std_logic ;
      MWRITEH_L       : IN     std_logic ;
      MWRITEL_L       : IN     std_logic ;
      PMDATAIN        : IN     LC3B_OWORD ;
      RESET_L         : IN     STD_LOGIC ;
      in_idlehit      : IN     std_logic ;
      in_load         : IN     std_logic ;
      in_writeback    : IN     std_logic ;
      DATAIN_internal : OUT    LC3b_word ;
      Dirty           : OUT    std_logic ;
      MRESP_H         : OUT    std_logic ;
      PMADDRESS       : OUT    LC3B_WORD ;
      PMDATAOUT       : OUT    LC3B_OWORD ;
      miss            : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Physical_Memory
   PORT (
      CLK       : IN     std_logic ;
      PMADDRESS : IN     LC3B_WORD ;
      PMDATAOUT : IN     LC3B_OWORD ;
      PMREAD_L  : IN     STD_LOGIC ;
      PMWRITE_L : IN     STD_LOGIC ;
      RESET_L   : IN     STD_LOGIC ;
      PMDATAIN  : OUT    LC3B_OWORD ;
      PMRESP_H  : OUT    STD_LOGIC 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Cache_Controller USE ENTITY ece411.Cache_Controller;
   FOR ALL : Cache_Datapath USE ENTITY ece411.Cache_Datapath;
   FOR ALL : Physical_Memory USE ENTITY ece411.Physical_Memory;
   -- pragma synthesis_on


BEGIN
   -- Architecture concurrent statements
   -- HDL Embedded Text Block 1 eb1
   MREAD_L <= instr_mread_l;
   MWRITEH_L <= '1';
   MWRITEL_L <= '1';
   Address <= instr_addr;
   instr_resp_h <= MRESP_H;
   
   instr_in <= DATAIN_internal;


   -- Instance port mappings.
   Cache_Cont : Cache_Controller
      PORT MAP (
         CLK          => CLK,
         Dirty        => Dirty,
         PMRESP_H     => PMRESP_H,
         RESET_L      => RESET_L,
         miss         => miss,
         PMREAD_L     => PMREAD_L,
         PMWRITE_L    => PMWRITE_L,
         in_idlehit   => in_idlehit,
         in_load      => in_load,
         in_writeback => in_writeback
      );
   Cache_DP1 : Cache_Datapath
      PORT MAP (
         Address         => Address,
         CLK             => CLK,
         Dataout         => Dataout,
         MREAD_L         => MREAD_L,
         MWRITEH_L       => MWRITEH_L,
         MWRITEL_L       => MWRITEL_L,
         PMDATAIN        => PMDATAIN,
         RESET_L         => RESET_L,
         in_idlehit      => in_idlehit,
         in_load         => in_load,
         in_writeback    => in_writeback,
         DATAIN_internal => DATAIN_internal,
         Dirty           => Dirty,
         MRESP_H         => MRESP_H,
         PMADDRESS       => PMADDRESS,
         PMDATAOUT       => PMDATAOUT,
         miss            => miss
      );
   PDRAM : Physical_Memory
      PORT MAP (
         CLK       => CLK,
         PMADDRESS => PMADDRESS,
         PMDATAOUT => PMDATAOUT,
         PMREAD_L  => PMREAD_L,
         PMWRITE_L => PMWRITE_L,
         RESET_L   => RESET_L,
         PMDATAIN  => PMDATAIN,
         PMRESP_H  => PMRESP_H
      );

END struct;
