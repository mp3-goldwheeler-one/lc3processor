configuration IR_config of IR is
   for untitled
   end for;
end IR_config;