configuration NZP_config of NZP is
   for untitled
   end for;
end NZP_config;